.title BGR Supply Sweep

*Libraries used
.lib $PDK_ROOT\/ihp-sg13g2/libs.tech/ngspice/models/cornerHBT.lib hbt_typ
.lib $PDK_ROOT\/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
.lib $PDK_ROOT\/ihp-sg13g2/libs.tech/ngspice/models/cornerRES.lib res_typ
.include ./bgr.cir.out

*Parameters 
.param resL=0.6u

*Ciruit under test
xbgr1 vdd vbg gnd bgr

*Supply 
V1 vdd gnd 1.3

*Temperature
.temp 27

*Analysis type
.dc V1 0 2.5 0.1

*Control statements
.control
run
cd simulationPlots
set hcopydevtype=svg
set color0=white
set color1=grey
set color2=red
hardcopy bgr_supply_sweep.svg v(vbg) title 'BGR Supply Sweep' ylabel 'Bandgap Reference Voltage' xlabel 'Supply Sweep' 
destroy all
quit
.endc
.end
